`ifndef DEFS_VH
`define DEFS_VH

// Field widths
`define INST_ID_W    16
`define SIZE_W       16
`define PRICE_W      32
`define TS_W         64

// Default configuration values
`define DEFAULT_IMB_THRESH       1
`define DEFAULT_MOMENTUM_DELTA   0
`define DEFAULT_MAX_SPREAD       1
`define DEFAULT_QTY              1
`define DEFAULT_MAX_POSITION     1000
`define DEFAULT_NOTIONAL_LIMIT   32'hFFFFFFFF

`endif // DEFS_VH
